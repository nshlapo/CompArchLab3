module testMem;
  initial begin
    $display("Testing memory");
  end
endmodule
